module topoclustering(clk, rst, io, eta, phi, et, e, eout, etout);
endmodule
